-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION Next_State_Logic_struct_config OF Next_State_Logic IS
   FOR struct
   END FOR;
END Next_State_Logic_struct_config;
