-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION my_xor_struct_config OF my_xor IS
   FOR struct
   END FOR;
END my_xor_struct_config;
