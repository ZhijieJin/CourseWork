-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION Vending_Machine_NAND_struct_config OF Vending_Machine_NAND IS
   FOR struct
   END FOR;
END Vending_Machine_NAND_struct_config;
