-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION Vending_Machine_struct_config OF Vending_Machine IS
   FOR struct
   END FOR;
END Vending_Machine_struct_config;
