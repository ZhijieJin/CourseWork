-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION Control_Logic_struct_config OF Control_Logic IS
   FOR struct
   END FOR;
END Control_Logic_struct_config;
